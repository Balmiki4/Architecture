module NotGate(input wire A, output wire o);

    assign o = ~A;

endmodule